error<=Linear_Audio xor Linear_Out;
